
module addertree_stage1(x14, x13, x12, x11, x10, x9, x8, x7, x6, x5, x4, x3, x2, x1, x0, 
                            );

input[8:0] x14, x13;
input[17:0] x12, x11;
input[35:0] x10, x9, x8, x7;
input[44:0] x6;
input[26:0] x5;
input[35:0] x4;
input[17:0] x3;
input[26:0] x2;
input[8:0] x1;
input[17:0] x0;

output o18, o17;
output [1:0] o16;
output [4:0] o15, o14;
output [6:0] o13;
output [8:0] o12;
output [9:0] o11;
output [10:0] o10;
output [11:0] o9;
output [10:0] o8;
output [9:0] o7;
output [9:0] o6;
output [8:0] o5;
output [7:0] o4;
output [5:0] o3;