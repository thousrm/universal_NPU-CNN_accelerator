
module adder_final(i19, i18, i17, i16, i15, i14, i13, i12, i11, i10, i9, i8, i7, i6, i5,
                    out);


input [1:0] i19, i18, i17, i16, i15, i14, i13, i12, i11, i10, i9, i8, i7, i6;
input i5;

wire [19:0] outb;

assign outb = (i19[0]<<19) + (i18[0]<<18) +(i17[0]<<17) +(i16[0]<<16) +(i15[0]<<15) +
                    (i14[0]<<14) +(i13[0]<<13) +(i12[0]<<12) +(i11[0]<<11) +
                    (i10[0]<<10) +(i9[0]<<9) +(i8[0]<<8) +(i7[0]<<7) +
                    (i6[0]<<6) +(i5<<5) + 
            (i19[1]<<19) + (i18[1]<<18) +(i17[1]<<17) +(i16[1]<<16) +(i15[1]<<15) +
                    (i14[1]<<14) +(i13[1]<<13) +(i12[1]<<12) +(i11[1]<<11) +
                    (i10[1]<<10) +(i9[1]<<9) +(i8[1]<<8) +(i7[1]<<7) +
                    (i6[1]<<6);


output [13:0] out;

assign out = outb[19-:14];

endmodule