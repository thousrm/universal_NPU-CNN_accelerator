
module _2cg(in, out);

input [7:0] in;
output [7:0] out;





endmodule