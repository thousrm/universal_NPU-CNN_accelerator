
module control_part();



endmodule