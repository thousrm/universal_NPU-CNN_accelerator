///////
//// - tx_top
//// - mac_lane
module mac (
    input logic
);



endmodule