///////
//// - tx_top
//// - mac_lane
module mac 
import tx_pkg::*;
(
    input logic
        
)
::



endmodule